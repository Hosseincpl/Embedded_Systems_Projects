-- RX and TX design
