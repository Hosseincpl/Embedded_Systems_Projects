-- 4 state parking lot
